LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUMADOR IS 
PORT 
(
SUMAX : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 );
SUMAY : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 );
CARRY_INS : IN STD_LOGIC;
CARRY_OUTS : BUFFER STD_LOGIC;
SUMA_sALIDA : OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0)
);
END SUMADOR;

ARCHITECTURE ARQUITECTURA_SUMA OF SUMADOR IS

--DECLARACION DE COMPONENTES -> SUMADOR UN BIT

COMPONENT SUMADOR_UN_BIT IS 
PORT 
(
A, B, CARRY_IN : IN STD_LOGIC;
SUM, CARRY_OUT : OUT STD_LOGIC
);
END COMPONENT;

SIGNAL C1 : STD_LOGIC;
SIGNAL C2 : STD_LOGIC;
SIGNAL C3 : STD_LOGIC;
SIGNAL C4 : STD_LOGIC;

BEGIN

SUMA1: SUMADOR_UN_BIT PORT MAP (A => SUMAX(0), B => SUMAY(0), CARRY_IN => CARRY_INS , SUM => SUMA_SALIDA(0), CARRY_OUT => C1);
SUMA2: SUMADOR_UN_BIT PORT MAP (A => SUMAX(1), B => SUMAY(1), CARRY_IN => C1 , SUM => SUMA_SALIDA(1), CARRY_OUT => C2);
SUMA3: SUMADOR_UN_BIT PORT MAP (A => SUMAX(2), B => SUMAY(2), CARRY_IN => C2 , SUM => SUMA_SALIDA(2), CARRY_OUT => C3);
SUMA4: SUMADOR_UN_BIT PORT MAP (A => SUMAX(3), B => SUMAY(3), CARRY_IN => C3 , SUM => SUMA_SALIDA(3), CARRY_OUT => CARRY_OUTS);

END ARQUITECTURA_SUMA;