LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUMADOR_UN_BIT IS 
PORT 
(
A, B, CARRY_IN : IN STD_LOGIC;
SUM, CARRY_OUT : OUT STD_LOGIC
);
END SUMADOR_UN_BIT;

ARCHITECTURE SUMADOR_UN_BIT OF SUMADOR_UN_BIT IS 
SIGNAL S1 : STD_LOGIC;
BEGIN 

S1 <= A XOR B;

SUM <= CARRY_IN XOR S1;

CARRY_OUT <= (CARRY_IN AND S1) OR ( A AND B);

END SUMADOR_UN_BIT;